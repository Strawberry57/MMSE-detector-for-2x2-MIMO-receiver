module qr_tb ();
   reg clk;
   reg reset;
   reg start;
   reg signed [15:0] h11,h12,h13,h14,h21,h22,h23,h24,h31,h32,h33,h34,h41,h42,h43,h44;

   wire signed [15:0] q11,q12,q13,q14,q21,q22,q23,q24,q31,q32,q33,q34,q41,q42,q43,q44,r11,r12,r13,r14,r22,r23,r24,r33,r34,r44;

   wire finish;

   qr qr(
      .clk (clk),
      .start (start),
      .reset (reset),
      .h11 (h11),
      .h12 (h12),
      .h13 (h13),
      .h14 (h14),
      .h21 (h21),
      .h22 (h22),
      .h23 (h23),
      .h24 (h24),
      .h31(h31),
      .h32 (h32),
      .h33 (h33),
      .h34 (h34),
      .h41 (h41),
      .h42 (h42),
      .h43 (h43),
      .h44 (h44),
      .q11 (q11),
      .q12 (q12),
      .q13 (q13),
      .q14 (q14),
      .q21 (q21),
      .q22 (q22),
      .q23 (q23),
      .q24 (q24),
      .q31 (q31),
      .q32 (q32),
      .q33 (q33),
      .q34 (q34),
      .q41 (q41),
      .q42 (q42),
      .q43 (q43),
      .q44 (q44),
      .r11 (r11),
      .r12 (r12),
      .r13 (r13),
      .r14 (r14),
      .r22 (r22),
      .r23 (r23),
      .r24 (r24),
      .r33 (r33),
      .r34 (r34),
      .r44 (r44),
      .q_a (q_a),
      .finish (finish)
   );

   initial begin
      reset = 1;
      #5 reset = 0;
      #10 reset = 1;
  end

   initial begin
      clk = 0;
      forever clk = #5 ~clk;
   end

   initial begin
      start = 1;
      h11 = 16'b00000010_00000000;
      h12 = 16'b00000001_00000000;
      h13 = 16'b00000010_00000000;
      h14 = 16'b00000001_00000000;
      h21 = 16'b00000001_00000000;
      h22 = 16'b00000010_00000000;
      h23 = 16'b00000001_00000000;
      h24 = 16'b00000010_00000000;
      h31 = 16'b00000101_00000000;
      h32 = 16'b00000001_00000000;
      h33 = 16'b00000011_00000000;
      h34 = 16'b00000001_00000000;
      h41 = 16'b00000011_00000000;
      h42 = 16'b00000101_00000000;
      h43 = 16'b00000001_00000000;
      h44 = 16'b00000011_00000000;
   
   end


endmodule